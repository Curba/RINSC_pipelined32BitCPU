// This is a common constants file for SystemVerilog macros to support the development
// in  Computer Architecture / Organization courses at METU Northern Cyprus Campus.
// Ali Muhtaroglu
// 

//////////////////////////////////////////
//              Constants               //
//////////////////////////////////////////

`define ON              1'b1
`define OFF             1'b0
`define ZERO            32'b0

